module tb();

initial begin

  run_test("test1");

end

endmodule
