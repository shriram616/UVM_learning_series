import uvm_pkg::*
`include "uvm_macros.svh";

`include "./top.sv"

//Test files
`include "../test/test1.sv"
  
 

