import uvm_pkg::*
`include "uvm_macros.svh";
package pkg;

  `include "./top.sv"

  //Test files
  `include "../test/test1.sv"
  
 
endpackage
